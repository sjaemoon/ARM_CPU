module mem_staged();