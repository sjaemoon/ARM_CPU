module branch_accel(clk, opcode, flag_wr_en, BrTaken, UncondBr, pc_rd)